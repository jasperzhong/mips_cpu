`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/06/03 01:12:15
// Design Name: 
// Module Name: CLZ
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CLZ(
    input [31:0] clz_in,
    output [31:0] clz_out
    );
    
    assign clz_out = 
        clz_in[31:31] == 1'b1 ? 32'd0:
        clz_in[31:30] == 2'b01 ? 32'd1:
        clz_in[31:29] == 3'b001 ? 32'd2:
        clz_in[31:28] == 4'b0001 ? 32'd3:
        clz_in[31:27] == 5'b00001 ? 32'd4:
        clz_in[31:26] == 6'b000001 ? 32'd5:
        clz_in[31:25] == 7'b0000001 ? 32'd6:
        clz_in[31:24] == 8'b00000001 ? 32'd7:
        clz_in[31:23] == 9'b000000001 ? 32'd8:
        clz_in[31:22] == 10'b0000000001 ? 32'd9:
        clz_in[31:21] == 11'b00000000001 ? 32'd10:
        clz_in[31:20] == 12'b000000000001 ? 32'd11:
        clz_in[31:19] == 13'b0000000000001 ? 32'd12:
        clz_in[31:18] == 14'b00000000000001 ? 32'd13:
        clz_in[31:17] == 15'b000000000000001 ? 32'd14:
        clz_in[31:16] == 16'b0000000000000001 ? 32'd15:
        clz_in[31:15] == 17'b00000000000000001 ? 32'd16:
        clz_in[31:14] == 18'b000000000000000001 ? 32'd17:
        clz_in[31:13] == 19'b0000000000000000001 ? 32'd18:
        clz_in[31:12] == 20'b00000000000000000001 ? 32'd19:
        clz_in[31:11] == 21'b000000000000000000001 ? 32'd20:
        clz_in[31:10] == 22'b0000000000000000000001 ? 32'd21:
        clz_in[31:9] == 23'b00000000000000000000001 ? 32'd22:
        clz_in[31:8] == 24'b000000000000000000000001 ? 32'd23:
        clz_in[31:7] == 25'b0000000000000000000000001 ? 32'd24:
        clz_in[31:6] == 26'b00000000000000000000000001 ? 32'd25:
        clz_in[31:5] == 27'b000000000000000000000000001 ? 32'd26:
        clz_in[31:4] == 28'b0000000000000000000000000001 ? 32'd27:
        clz_in[31:3] == 29'b00000000000000000000000000001 ? 32'd28:
        clz_in[31:2] == 30'b000000000000000000000000000001 ? 32'd29:
        clz_in[31:1] == 31'b0000000000000000000000000000001 ? 32'd30:
        clz_in[31:0] == 32'b00000000000000000000000000000001 ? 32'd31:
        32'd32;
endmodule
